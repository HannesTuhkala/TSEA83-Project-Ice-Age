library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity cpu is
	port (
		clk: in std_logic;
		a1 : in ???;
		a2 : out ???);
end cpu;

architecture behavioral of cpu is
	
	----------------------------------------------------
	---------------------PROGRAM_MEMORY-----------------
	----------------------------------------------------
	-- Declaration of a doubleported block-RAM
	-- with 512 addresses of 32 bits width.
	type pm_t is array(0 to 511) of
		std_logic_vector(31 downto 0);
		
	-- Reset all bits on all adresses
	signal pm : pm_t := (others => (others => '0'));
	
	-- port 1
	signal adress1 : std_logic_vector(8 downto 0);
	signal rw1 : std_logic; -- Read/Write flag for port 1
	signal ce1 : std_logic; -- Count enable flag for port 1
	signal data1 : std_logic_vector(31 downto 0); -- Our instruction, which is 32 bits long.
	
	-- port 2
	signal adress2 : std_logic_vector(8 downto 0);
	signal rw2 : std_logic; -- Read/Write flag for port 2
	signal ce2 : std_logic; -- Count enable flag for port 2
	signal data2 : std_logic_vector(31 downto 0)); -- Our instruction, which is 32 bits long.

	--------------------------------------------------
	--------------END OF PROGRAM MEMORY---------------
	--------------------------------------------------

begin

	-------- Program Memory ---------
	PROCESS(clk)
	BEGIN
		if (rising_edge(clk)) then
			if (re1 = '0') then
				data1 <= (adress1);
			end if;
		end if;
	END PROCESS;
	-------- END Program Memory -------


end behavioral;
