entity graphic
	port (
		b1 : in ???;
		b2 : out ???;
		b3 : out ???);
end graphic;

architecture behavioral of graphic is

begin

end behavioral;