entity cpu
	port (
		a1 : in ???
		a2 : out ???);
end CPU;

architecture behavioral of cpu is

begin

end behavioral;